import FIFO::*;