// This file contains types used in the compression function

// Control Word types



typedef Bit#(6) ShiftFactor;